module basic_control(

);

endmodule
