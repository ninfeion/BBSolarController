// Verilog created by ORCAD Capture

module EP4CE6E144 
 ( 
 );


initial
	begin
	end

endmodule
